module signExtend(
  input [31:0] immSel,
  input [31:0] in, // todo: 20 ig
  output [31:0] out
);
endmodule